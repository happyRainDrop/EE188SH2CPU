--Hello
--
--This is Nerissa's personal log